module playingcards

import rand
